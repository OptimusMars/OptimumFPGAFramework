package helper_func;
  


  
endpackage : helper_func