// Static clock divisor
module clkdiv_s #(parameter DIVISOR = 3) (
  input  clk ,
  input  rst ,
  output clko
);

endmodule