package mult_pkg;

function integer rtoi (input integer x);
  rtoi = x;
endfunction

function longint pow2repr(real value);
  


endfunction

  

endpackage : mult_pkg

